module groblon_core


import os
import time





pub fn file_watcher()
{
  // Todo
}