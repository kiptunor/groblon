module config_utils



struct Config
{
  // Config fields soon
}

pub fn load_config()
{
  // Load and return config structure
}

pub fn save_config(config: Config)
{
  // Save config structure to file
}
