module main


import server_api
import groblon_utils



fn main()
{
  server_api.server_init()
  // println(groblon_utils.get_default_note_dir())
  // println(groblon_utils.get_config_dir())
  
  // groblon_utils.setup()
}
