module main


import server_api



fn main()
{
  server_api.server_init()
}
