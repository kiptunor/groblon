module main



import groblon_core



fn main()
{
  groblon_core.setup()
  
  server_init()
}
